-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
--                                                                           --
-- File Name: TB_Network_Detection.vhd                                                  --
-- Author: Phillip Jones (phjones@iastate.edu  )                             --
-- Date: 2/1/2018                                                           --
--                                                                           --
-- Description: Base testbench for generating stimulus input for             -- 
-- DUT  (Device Under Test)                                                  --
--                                                                           --
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity ppm_tb_gen is
port
(
my_in : in std_logic -- input needed to keep modelsim from complainning???
);
end ppm_tb_gen;

architecture tb1 of ppm_tb_gen is

----------------------------------------------
--       Component declarations             --
----------------------------------------------

-- Device under test

component ppm_generation is
	port (
		-- Users to add ports here
        	PPM_OUT  : out std_logic;
        	PPM_CLK  : in std_logic;
		S_AXI_ARESETN : in std_logic;
		slv_reg0 : in std_logic_vector(31 downto 0);
		slv_reg10 : in std_logic_vector(31 downto 0);
		slv_reg11 : in std_logic_vector(31 downto 0);
		slv_reg12 : in std_logic_vector(31 downto 0);
		slv_reg13 : in std_logic_vector(31 downto 0);
		slv_reg14 : in std_logic_vector(31 downto 0);
		slv_reg15 : in std_logic_vector(31 downto 0)
	);
end component ppm_generation;



----------------------------------------------
--          Signal declarations             --
----------------------------------------------
type my_input_states is (S0, S1, S2, S3, S4, S5, S6, S7, S8, S9, S10, S11, 
                         S12, S13, S14, S15, S16, S17, S18, S19, S20, S21, 
			S22,S23,S24,S25,S26,S27,S28,S29, STOP_TEST);

	signal ppm : std_logic;
	signal reset : std_logic;
	signal clk : std_logic;
	signal input_state    : my_input_states;  -- Direct which input vector to use



begin


-- Processes


------------------------------------------------------------
------------------------------------------------------------
--                                                        --
-- Process Name: DUT stimulus                             --
--                                                        --
-- Send inputs to dut. Holds inputs for HOLD_INPUT_reg    --
--  clk cycles                                            --
--                                                        --
------------------------------------------------------------
------------------------------------------------------------
ppm_stimulus : process(clk)
begin
  if (clk = '1' and clk'event) then

    -- Initialize the test
    if(reset = '0') then
      --input_state    <= S0;
    end if;
	
	case input_state is
		when S0 => 
			reset <= '0';
			input_state <= S1;
		when S1 =>
			reset <= '1';
			input_state <= S2;
		when S2 => 

		when others =>
	end case;
  end if;
end process ppm_stimulus;



-- Combinational assignments

  -- none

-- Connect DUT (Network Detection circuit) to the testbench

my_ppm_gen : ppm_generation
port map
(
        	PPM_OUT  => ppm,
        	PPM_CLK  => clk,
		S_AXI_ARESETN => reset,
		slv_reg0 => x"00000000",
		--slv_reg10 => x"000186A0",
		slv_reg10 => x"00000004",
		slv_reg11 => x"00000004",
		slv_reg12 => x"00000004",
		slv_reg13 => x"00000004",
		slv_reg14 => x"00000004",
		slv_reg15 => x"00000004"
);


end tb1;
